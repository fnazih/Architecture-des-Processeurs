-------------------------------------------------------------------------------
-- Title      : DLX_top
-- Project    : 
-------------------------------------------------------------------------------
-- File       : DLX_top.vhd
-- Author     :   <michel agoyan@ROU13572>
-- Company    : 
-- Created    : 2015-11-25
-- Last update: 2019-12-03
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: DLX data path + control path
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2015-11-25  1.0      michel agoyan   Created
-- 2019-08-21  1.1      Olivier potin   Modified to implement RISCV Monocycle
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use work.RV32I_components.all;

entity RV32I_Monocycle_top is

  port (
    clk_i    : in std_logic;
    resetn_i : in std_logic);

end entity RV32I_Monocycle_top;

architecture RV32I_Monocycle_top_architecture of RV32I_Monocycle_top is
  
-- RV32 current instruction (i.e from datapath to control path) 
-- see Patterson & Hennessy page  257 for global sheme
  signal Instruction_s : std_logic_vector(31 downto 0);

  
-- outputs signal generated by controler (i.e from controlpath to datapath)
-- see patterson and Hennessy page 256
 
  signal alu_control_s : std_logic_vector(3 downto 0);
  signal reg_write_s   : std_logic;
  signal alu_src1_s    : std_logic_vector(1 downto 0);
  signal alu_src2_s    : std_logic_vector(0 downto 0);
  signal imm_gen_sel_s : std_logic_vector(1 downto 0);
  signal alu_zero_s   : std_logic;
  signal alu_lt_s      : std_logic;
 
  
begin  -- architecture RV32I_Monocycle_top_architecture

  RV32I_Monocycle_controlpath_1: RV32I_Monocycle_controlpath
    port map (
      instruction_i => instruction_s,
      alu_zero_i    => alu_zero_s,
      alu_lt_i      => alu_lt_s,
      alu_src1_o    => alu_src1_s,
      alu_src2_o    => alu_src2_s,
      alu_control_o => alu_control_s,
      imm_gen_sel_o => imm_gen_sel_s,
      reg_write_o   => reg_write_s);

  RV32I_Monocycle_datapath_1 : RV32I_Monocycle_datapath
    port map (
      clk_i         => clk_i,
      resetn_i      => resetn_i,
      alu_control_i => alu_control_s,
      reg_write_i   => reg_write_s,
      alu_src1_i    => alu_src1_s,
      alu_src2_i    => alu_src2_s,
      imm_gen_sel_i => imm_gen_sel_s,
      instruction_o => instruction_s,
      alu_zero_o    => alu_zero_s,
      alu_lt_o      => alu_lt_s);
end architecture RV32I_Monocycle_top_architecture;
